`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Assignment 6
// Group 69
// Team Member 1: Rushil Venkateswar (20CS30045)
// Team Member 2: Jatin Gupta (20CS10087)
// SEM 5 (Autumn 2022-23)
//////////////////////////////////////////////////////////////////////////////////

module diff_module(input [31:0] in, output [31:0] out);
    always @(*) begin
        case(in)
            32'b00000000000000000000000000000000: out = 32'b00000000000000000000000000100001;
            32'b00000000000000000000000000000001: out = 32'b00000000000000000000000000000001;
            32'b00000000000000000000000000000010: out = 32'b00000000000000000000000000000010;
            32'b00000000000000000000000000000100: out = 32'b00000000000000000000000000000011;
            32'b00000000000000000000000000001000: out = 32'b00000000000000000000000000000100;
            32'b00000000000000000000000000010000: out = 32'b00000000000000000000000000000101;
            32'b00000000000000000000000000100000: out = 32'b00000000000000000000000000000110;
            32'b00000000000000000000000001000000: out = 32'b00000000000000000000000000000111;
            32'b00000000000000000000000010000000: out = 32'b00000000000000000000000000001000;
            32'b00000000000000000000000100000000: out = 32'b00000000000000000000000000001001;
            32'b00000000000000000000001000000000: out = 32'b00000000000000000000000000001010;
            32'b00000000000000000000010000000000: out = 32'b00000000000000000000000000001011;
            32'b00000000000000000000100000000000: out = 32'b00000000000000000000000000001100;
            32'b00000000000000000001000000000000: out = 32'b00000000000000000000000000001101;
            32'b00000000000000000010000000000000: out = 32'b00000000000000000000000000001110;
            32'b00000000000000000100000000000000: out = 32'b00000000000000000000000000001111;
            32'b00000000000000001000000000000000: out = 32'b00000000000000000000000000010000;
            32'b00000000000000010000000000000000: out = 32'b00000000000000000000000000010001;
            32'b00000000000000100000000000000000: out = 32'b00000000000000000000000000010010;
            32'b00000000000001000000000000000000: out = 32'b00000000000000000000000000010011;
            32'b00000000000010000000000000000000: out = 32'b00000000000000000000000000010100;
            32'b00000000000100000000000000000000: out = 32'b00000000000000000000000000010101;
            32'b00000000001000000000000000000000: out = 32'b00000000000000000000000000010110;
            32'b00000000010000000000000000000000: out = 32'b00000000000000000000000000010111;
            32'b00000000100000000000000000000000: out = 32'b00000000000000000000000000011000;
            32'b00000001000000000000000000000000: out = 32'b00000000000000000000000000011001;
            32'b00000010000000000000000000000000: out = 32'b00000000000000000000000000011010;
            32'b00000100000000000000000000000000: out = 32'b00000000000000000000000000011011;
            32'b00001000000000000000000000000000: out = 32'b00000000000000000000000000011100;
            32'b00010000000000000000000000000000: out = 32'b00000000000000000000000000011101;
            32'b00100000000000000000000000000000: out = 32'b00000000000000000000000000011110;
            32'b01000000000000000000000000000000: out = 32'b00000000000000000000000000011111;
            32'b10000000000000000000000000000000: out = 32'b00000000000000000000000000100000;
        endcase
    end
endmodule
            

            