`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Assignment 6
// Group 69
// Team Member 1: Rushil Venkateswar (20CS30045)
// Team Member 2: Jatin Gupta (20CS10087)
// SEM 5 (Autumn 2022-23)
//////////////////////////////////////////////////////////////////////////////////

module diff_module(input [31:0] in, output reg [31:0] out);
    always @(*) begin
        case(in)
            32'b00000000000000000000000000000000:begin out = 32'b00000000000000000000000000000000; end
            32'b00000000000000000000000000000001:begin out = 32'b00000000000000000000000000000001; end
            32'b00000000000000000000000000000010:begin out = 32'b00000000000000000000000000000010; end
            32'b00000000000000000000000000000100:begin out = 32'b00000000000000000000000000000011; end
            32'b00000000000000000000000000001000:begin out = 32'b00000000000000000000000000000100; end
            32'b00000000000000000000000000010000:begin out = 32'b00000000000000000000000000000101; end
            32'b00000000000000000000000000100000:begin out = 32'b00000000000000000000000000000110; end
            32'b00000000000000000000000001000000:begin out = 32'b00000000000000000000000000000111; end
            32'b00000000000000000000000010000000:begin out = 32'b00000000000000000000000000001000; end
            32'b00000000000000000000000100000000:begin out = 32'b00000000000000000000000000001001; end
            32'b00000000000000000000001000000000:begin out = 32'b00000000000000000000000000001010; end
            32'b00000000000000000000010000000000:begin out = 32'b00000000000000000000000000001011; end
            32'b00000000000000000000100000000000:begin out = 32'b00000000000000000000000000001100; end
            32'b00000000000000000001000000000000:begin out = 32'b00000000000000000000000000001101; end
            32'b00000000000000000010000000000000:begin out = 32'b00000000000000000000000000001110; end
            32'b00000000000000000100000000000000:begin out = 32'b00000000000000000000000000001111; end
            32'b00000000000000001000000000000000:begin out = 32'b00000000000000000000000000010000; end
            32'b00000000000000010000000000000000:begin out = 32'b00000000000000000000000000010001; end
            32'b00000000000000100000000000000000:begin out = 32'b00000000000000000000000000010010; end
            32'b00000000000001000000000000000000:begin out = 32'b00000000000000000000000000010011; end
            32'b00000000000010000000000000000000:begin out = 32'b00000000000000000000000000010100; end
            32'b00000000000100000000000000000000:begin out = 32'b00000000000000000000000000010101; end
            32'b00000000001000000000000000000000:begin out = 32'b00000000000000000000000000010110; end
            32'b00000000010000000000000000000000:begin out = 32'b00000000000000000000000000010111; end
            32'b00000000100000000000000000000000:begin out = 32'b00000000000000000000000000011000; end
            32'b00000001000000000000000000000000:begin out = 32'b00000000000000000000000000011001; end
            32'b00000010000000000000000000000000:begin out = 32'b00000000000000000000000000011010; end
            32'b00000100000000000000000000000000:begin out = 32'b00000000000000000000000000011011; end
            32'b00001000000000000000000000000000:begin out = 32'b00000000000000000000000000011100; end
            32'b00010000000000000000000000000000:begin out = 32'b00000000000000000000000000011101; end
            32'b00100000000000000000000000000000:begin out = 32'b00000000000000000000000000011110; end
            32'b01000000000000000000000000000000:begin out = 32'b00000000000000000000000000011111; end
            32'b10000000000000000000000000000000:begin out = 32'b00000000000000000000000000100000; end
				default: out = 32'b0;
        endcase
    end
endmodule
        