module dff_structural(input [3:0] set, input [3:0] Clk, input [3:0] Data, output  )